** Profile: "SCHEMATIC1-Time-domain-sim"  [ C:\USERS\BENJAMIN BEAUDOIN\DOCUMENTS\GITHUB\ALTIUM-GITHUB-REPO-BEAUD082\ALTIUM PROJECTS FILES\ORCAD_SIM_FILES\independent study simulation test-pspicefiles\schematic1\time-domain-sim.sim ] 

** Creating circuit file "Time-domain-sim.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
* From [PSPICE NETLIST] section of C:\SPB_Data\cdssetup\OrCAD_PSpice/16.6.0/PSpice.ini file:
.lib "nomd.lib" 

*Analysis directives: 
.TRAN  0 100us 0 
.OPTIONS ADVCONV
.PROBE64 V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\SCHEMATIC1.net" 


.END
